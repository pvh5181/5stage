module Counter4bit_Up(
	input clk_50M,
	input load,
	input enable,
	output [6:0] display
);

reg [3:0] out_CNT;
wire clk_1;
wire load_new;
always @(posedge clk_1)
begin
	if(enable)
		if(load_new)
			out_CNT = 0;
		else
			begin
				out_CNT <= out_CNT +1;
			end

end


clock_divider(clk_50M, clk_1);
edge_detection(clk_50M, clk_1, load, load_new);
seven_segment_display a(out_CNT[3:0], display);

endmodule